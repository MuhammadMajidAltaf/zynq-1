---------------------------------------------------------------------------
-- Author   : Ali Lown <ali@lown.me.uk>
-- File          : offload_top.vhdl
--
-- Abstract :
--
---------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.all;

---------------------------------------------------------------------------
Entity offload_top is 
---------------------------------------------------------------------------
port 
(
  clk : in std_logic;
  reset_n : in std_logic;

  s_axis_tvalid : in std_logic;
  s_axis_tready : out std_logic;
  s_axis_tdata : in std_logic_vector(31 downto 0);
  s_axis_tkeep : in std_logic_vector(3 downto 0);
  s_axis_tlast : in std_logic;

  m_axis_tvalid : out std_logic;
  m_axis_tready : in std_logic;
  m_axis_tdata : out std_logic_vector(31 downto 0);
  m_axis_tkeep : out std_logic_vector(3 downto 0);
  m_axis_tlast : out std_logic;
  dbg : out std_logic_vector(3 downto 0)
);
end entity;


---------------------------------------------------------------------------
Architecture offload_top_1 of offload_top is
---------------------------------------------------------------------------

  type state_type is (s0_check, s1_have_header, s2_compute, s3_results);
  signal state : state_type;

  --ignoring SP, LR, PC registers
  type reg_array is array (0 to 13) of std_logic_vector(31 downto 0);
  signal regs_in, regs_out : reg_array;
  signal reg_count : natural := 0;
  signal s_axis_tready_out : std_logic;

  constant PKT_MAGIC : std_logic_vector(31 downto 0) := x"0FFA0FFB";

--<<< BEGIN SIGNALS
signal t_40_s, t_50_s, t_60_s, t_70_s, t_80_s, t_90_s, t_a0_s, t_b0_s, t_c0_s, t_d0_s, r0_dc, r1_dc, r2_dc, r3_dc, r4_dc, r5_dc, r6_dc, r7_dc, r8_dc, r9_dc, r10_dc, r11_dc, r12_dc, r13_dc, r0_3c, r1_3c, r2_3c, r3_3c, r4_3c, r5_3c, r6_3c, r7_3c, r8_3c, r9_3c, r10_3c, r11_3c, r12_3c, r13_3c, r0_40, r1_40, r2_40, r3_40, r4_40, r5_40, r6_40, r7_40, r8_40, r9_40, r10_40, r11_40, r12_40, r13_40, r0_44, r1_44, r2_44, r3_44, r4_44, r5_44, r6_44, r7_44, r8_44, r9_44, r10_44, r11_44, r12_44, r13_44, r0_48, r1_48, r2_48, r3_48, r4_48, r5_48, r6_48, r7_48, r8_48, r9_48, r10_48, r11_48, r12_48, r13_48, r0_4c, r1_4c, r2_4c, r3_4c, r4_4c, r5_4c, r6_4c, r7_4c, r8_4c, r9_4c, r10_4c, r11_4c, r12_4c, r13_4c, r0_50, r1_50, r2_50, r3_50, r4_50, r5_50, r6_50, r7_50, r8_50, r9_50, r10_50, r11_50, r12_50, r13_50, r0_54, r1_54, r2_54, r3_54, r4_54, r5_54, r6_54, r7_54, r8_54, r9_54, r10_54, r11_54, r12_54, r13_54, r0_58, r1_58, r2_58, r3_58, r4_58, r5_58, r6_58, r7_58, r8_58, r9_58, r10_58, r11_58, r12_58, r13_58, r0_5c, r1_5c, r2_5c, r3_5c, r4_5c, r5_5c, r6_5c, r7_5c, r8_5c, r9_5c, r10_5c, r11_5c, r12_5c, r13_5c, r0_60, r1_60, r2_60, r3_60, r4_60, r5_60, r6_60, r7_60, r8_60, r9_60, r10_60, r11_60, r12_60, r13_60, r0_64, r1_64, r2_64, r3_64, r4_64, r5_64, r6_64, r7_64, r8_64, r9_64, r10_64, r11_64, r12_64, r13_64, r0_68, r1_68, r2_68, r3_68, r4_68, r5_68, r6_68, r7_68, r8_68, r9_68, r10_68, r11_68, r12_68, r13_68, r0_6c, r1_6c, r2_6c, r3_6c, r4_6c, r5_6c, r6_6c, r7_6c, r8_6c, r9_6c, r10_6c, r11_6c, r12_6c, r13_6c, r0_70, r1_70, r2_70, r3_70, r4_70, r5_70, r6_70, r7_70, r8_70, r9_70, r10_70, r11_70, r12_70, r13_70, r0_74, r1_74, r2_74, r3_74, r4_74, r5_74, r6_74, r7_74, r8_74, r9_74, r10_74, r11_74, r12_74, r13_74, r0_78, r1_78, r2_78, r3_78, r4_78, r5_78, r6_78, r7_78, r8_78, r9_78, r10_78, r11_78, r12_78, r13_78, r0_7c, r1_7c, r2_7c, r3_7c, r4_7c, r5_7c, r6_7c, r7_7c, r8_7c, r9_7c, r10_7c, r11_7c, r12_7c, r13_7c, r0_80, r1_80, r2_80, r3_80, r4_80, r5_80, r6_80, r7_80, r8_80, r9_80, r10_80, r11_80, r12_80, r13_80, r0_84, r1_84, r2_84, r3_84, r4_84, r5_84, r6_84, r7_84, r8_84, r9_84, r10_84, r11_84, r12_84, r13_84, r0_88, r1_88, r2_88, r3_88, r4_88, r5_88, r6_88, r7_88, r8_88, r9_88, r10_88, r11_88, r12_88, r13_88, r0_8c, r1_8c, r2_8c, r3_8c, r4_8c, r5_8c, r6_8c, r7_8c, r8_8c, r9_8c, r10_8c, r11_8c, r12_8c, r13_8c, r0_90, r1_90, r2_90, r3_90, r4_90, r5_90, r6_90, r7_90, r8_90, r9_90, r10_90, r11_90, r12_90, r13_90, r0_94, r1_94, r2_94, r3_94, r4_94, r5_94, r6_94, r7_94, r8_94, r9_94, r10_94, r11_94, r12_94, r13_94, r0_98, r1_98, r2_98, r3_98, r4_98, r5_98, r6_98, r7_98, r8_98, r9_98, r10_98, r11_98, r12_98, r13_98, r0_9c, r1_9c, r2_9c, r3_9c, r4_9c, r5_9c, r6_9c, r7_9c, r8_9c, r9_9c, r10_9c, r11_9c, r12_9c, r13_9c, r0_a0, r1_a0, r2_a0, r3_a0, r4_a0, r5_a0, r6_a0, r7_a0, r8_a0, r9_a0, r10_a0, r11_a0, r12_a0, r13_a0, r0_a4, r1_a4, r2_a4, r3_a4, r4_a4, r5_a4, r6_a4, r7_a4, r8_a4, r9_a4, r10_a4, r11_a4, r12_a4, r13_a4, r0_a8, r1_a8, r2_a8, r3_a8, r4_a8, r5_a8, r6_a8, r7_a8, r8_a8, r9_a8, r10_a8, r11_a8, r12_a8, r13_a8, r0_ac, r1_ac, r2_ac, r3_ac, r4_ac, r5_ac, r6_ac, r7_ac, r8_ac, r9_ac, r10_ac, r11_ac, r12_ac, r13_ac, r0_b0, r1_b0, r2_b0, r3_b0, r4_b0, r5_b0, r6_b0, r7_b0, r8_b0, r9_b0, r10_b0, r11_b0, r12_b0, r13_b0, r0_b4, r1_b4, r2_b4, r3_b4, r4_b4, r5_b4, r6_b4, r7_b4, r8_b4, r9_b4, r10_b4, r11_b4, r12_b4, r13_b4, r0_b8, r1_b8, r2_b8, r3_b8, r4_b8, r5_b8, r6_b8, r7_b8, r8_b8, r9_b8, r10_b8, r11_b8, r12_b8, r13_b8, r0_bc, r1_bc, r2_bc, r3_bc, r4_bc, r5_bc, r6_bc, r7_bc, r8_bc, r9_bc, r10_bc, r11_bc, r12_bc, r13_bc, r0_c0, r1_c0, r2_c0, r3_c0, r4_c0, r5_c0, r6_c0, r7_c0, r8_c0, r9_c0, r10_c0, r11_c0, r12_c0, r13_c0, r0_c4, r1_c4, r2_c4, r3_c4, r4_c4, r5_c4, r6_c4, r7_c4, r8_c4, r9_c4, r10_c4, r11_c4, r12_c4, r13_c4, r0_c8, r1_c8, r2_c8, r3_c8, r4_c8, r5_c8, r6_c8, r7_c8, r8_c8, r9_c8, r10_c8, r11_c8, r12_c8, r13_c8, r0_cc, r1_cc, r2_cc, r3_cc, r4_cc, r5_cc, r6_cc, r7_cc, r8_cc, r9_cc, r10_cc, r11_cc, r12_cc, r13_cc, r0_d0, r1_d0, r2_d0, r3_d0, r4_d0, r5_d0, r6_d0, r7_d0, r8_d0, r9_d0, r10_d0, r11_d0, r12_d0, r13_d0, r0_d4, r1_d4, r2_d4, r3_d4, r4_d4, r5_d4, r6_d4, r7_d4, r8_d4, r9_d4, r10_d4, r11_d4, r12_d4, r13_d4, r0_d8, r1_d8, r2_d8, r3_d8, r4_d8, r5_d8, r6_d8, r7_d8, r8_d8, r9_d8, r10_d8, r11_d8, r12_d8, r13_d8 : std_logic_vector(31 downto 0);
--->>> END SIGNALS

begin

  s_axis_tready <= s_axis_tready_out;

  FSM: process(clk, reset_n, s_axis_tvalid, s_axis_tkeep, s_axis_tdata, m_axis_tready)
  begin
    if clk'event and clk='1' then
      if reset_n = '0' then
        state <= s0_check;
        s_axis_tready_out <= '0';
        m_axis_tvalid <= '0';
        reg_count <= 0;
        dbg <= "0000";
      else
        case state is
          when s0_check =>
            s_axis_tready_out <= '1';
            m_axis_tvalid <= '0';
            m_axis_tlast <= '0';

            if s_axis_tvalid = '1' then
              if s_axis_tkeep = "0000" and s_axis_tdata = PKT_MAGIC then
                reg_count <= 0;
                state <= s1_have_header;
              end if;
            end if;

          when s1_have_header =>
            dbg(1) <= '1';

            --Next 14 data items are the register starting states - assuming no partial packets
            if not (s_axis_tkeep = "1111" ) or s_axis_tlast = '1' or s_axis_tvalid = '0' then
              state <= s0_check;
            else
              regs_in(reg_count) <= s_axis_tdata;
              if reg_count = 13 then
                state <= s2_compute;
              else
                reg_count <= reg_count + 1;
              end if;
            end if;

          when s2_compute =>
            dbg(3) <= '1';
            state <= s3_results;
            reg_count <= 0;

          when s3_results =>
            m_axis_tvalid <= '1';
            m_axis_tkeep <= "1111";
            if m_axis_tready = '1' then
              m_axis_tlast <= '0';
              if reg_count = 0 then
                m_axis_tdata <= PKT_MAGIC;
              else
                m_axis_tdata <= regs_out(reg_count-1);
              end if;
              if reg_count = 14 then
                m_axis_tlast <= '1';
                state <= s0_check;
              else
                reg_count <= reg_count + 1;
              end if;
            end if;

        end case;
      end if;
    end if;
  end process;

---<<< BEGIN LOGIC
r0_3c <= regs_in(0);
r1_3c <= regs_in(1);
r2_3c <= regs_in(2);
r3_3c <= regs_in(3);
r4_3c <= regs_in(4);
r5_3c <= regs_in(5);
r6_3c <= regs_in(6);
r7_3c <= regs_in(7);
r8_3c <= regs_in(8);
r9_3c <= regs_in(9);
r10_3c <= regs_in(10);
r11_3c <= regs_in(11);
r12_3c <= regs_in(12);
r13_3c <= regs_in(13);
r3_40 <= std_logic_vector( unsigned(r0_3c) + unsigned(r1_3c));
r0_40 <= r0_3c;
r1_40 <= r1_3c;
r2_40 <= r2_3c;
r4_40 <= r4_3c;
r5_40 <= r5_3c;
r6_40 <= r6_3c;
r7_40 <= r7_3c;
r8_40 <= r8_3c;
r9_40 <= r9_3c;
r10_40 <= r10_3c;
r11_40 <= r11_3c;
r12_40 <= r12_3c;
r13_40 <= r13_3c;
t_40_s <= std_logic_vector(unsigned(r3_40) sll TO_INTEGER(unsigned(r0_40)));
r3_44 <= std_logic_vector( unsigned(r1_40) or unsigned(t_40_s));
r0_44 <= r0_40;
r1_44 <= r1_40;
r2_44 <= r2_40;
r4_44 <= r4_40;
r5_44 <= r5_40;
r6_44 <= r6_40;
r7_44 <= r7_40;
r8_44 <= r8_40;
r9_44 <= r9_40;
r10_44 <= r10_40;
r11_44 <= r11_40;
r12_44 <= r12_40;
r13_44 <= r13_40;
r3_48 <= std_logic_vector( unsigned(r3_44) xor unsigned(r0_44));
r0_48 <= r0_44;
r1_48 <= r1_44;
r2_48 <= r2_44;
r4_48 <= r4_44;
r5_48 <= r5_44;
r6_48 <= r6_44;
r7_48 <= r7_44;
r8_48 <= r8_44;
r9_48 <= r9_44;
r10_48 <= r10_44;
r11_48 <= r11_44;
r12_48 <= r12_44;
r13_48 <= r13_44;
r3_4c <= std_logic_vector( unsigned(r3_48) - unsigned(r1_48));
r0_4c <= r0_48;
r1_4c <= r1_48;
r2_4c <= r2_48;
r4_4c <= r4_48;
r5_4c <= r5_48;
r6_4c <= r6_48;
r7_4c <= r7_48;
r8_4c <= r8_48;
r9_4c <= r9_48;
r10_4c <= r10_48;
r11_4c <= r11_48;
r12_4c <= r12_48;
r13_4c <= r13_48;
r3_50 <= std_logic_vector(RESIZE(unsigned(r3_4c) * unsigned(r0_4c) + unsigned(r1_4c), 32));
r0_50 <= r0_4c;
r1_50 <= r1_4c;
r2_50 <= r2_4c;
r4_50 <= r4_4c;
r5_50 <= r5_4c;
r6_50 <= r6_4c;
r7_50 <= r7_4c;
r8_50 <= r8_4c;
r9_50 <= r9_4c;
r10_50 <= r10_4c;
r11_50 <= r11_4c;
r12_50 <= r12_4c;
r13_50 <= r13_4c;
t_50_s <= std_logic_vector(unsigned(r3_50) sll TO_INTEGER(unsigned(r0_50)));
r3_54 <= std_logic_vector( unsigned(r1_50) or unsigned(t_50_s));
r0_54 <= r0_50;
r1_54 <= r1_50;
r2_54 <= r2_50;
r4_54 <= r4_50;
r5_54 <= r5_50;
r6_54 <= r6_50;
r7_54 <= r7_50;
r8_54 <= r8_50;
r9_54 <= r9_50;
r10_54 <= r10_50;
r11_54 <= r11_50;
r12_54 <= r12_50;
r13_54 <= r13_50;
r3_58 <= std_logic_vector( unsigned(r3_54) xor unsigned(r0_54));
r0_58 <= r0_54;
r1_58 <= r1_54;
r2_58 <= r2_54;
r4_58 <= r4_54;
r5_58 <= r5_54;
r6_58 <= r6_54;
r7_58 <= r7_54;
r8_58 <= r8_54;
r9_58 <= r9_54;
r10_58 <= r10_54;
r11_58 <= r11_54;
r12_58 <= r12_54;
r13_58 <= r13_54;
r3_5c <= std_logic_vector( unsigned(r3_58) - unsigned(r1_58));
r0_5c <= r0_58;
r1_5c <= r1_58;
r2_5c <= r2_58;
r4_5c <= r4_58;
r5_5c <= r5_58;
r6_5c <= r6_58;
r7_5c <= r7_58;
r8_5c <= r8_58;
r9_5c <= r9_58;
r10_5c <= r10_58;
r11_5c <= r11_58;
r12_5c <= r12_58;
r13_5c <= r13_58;
r3_60 <= std_logic_vector(RESIZE(unsigned(r3_5c) * unsigned(r0_5c) + unsigned(r1_5c), 32));
r0_60 <= r0_5c;
r1_60 <= r1_5c;
r2_60 <= r2_5c;
r4_60 <= r4_5c;
r5_60 <= r5_5c;
r6_60 <= r6_5c;
r7_60 <= r7_5c;
r8_60 <= r8_5c;
r9_60 <= r9_5c;
r10_60 <= r10_5c;
r11_60 <= r11_5c;
r12_60 <= r12_5c;
r13_60 <= r13_5c;
t_60_s <= std_logic_vector(unsigned(r3_60) sll TO_INTEGER(unsigned(r0_60)));
r3_64 <= std_logic_vector( unsigned(r1_60) or unsigned(t_60_s));
r0_64 <= r0_60;
r1_64 <= r1_60;
r2_64 <= r2_60;
r4_64 <= r4_60;
r5_64 <= r5_60;
r6_64 <= r6_60;
r7_64 <= r7_60;
r8_64 <= r8_60;
r9_64 <= r9_60;
r10_64 <= r10_60;
r11_64 <= r11_60;
r12_64 <= r12_60;
r13_64 <= r13_60;
r3_68 <= std_logic_vector( unsigned(r3_64) xor unsigned(r0_64));
r0_68 <= r0_64;
r1_68 <= r1_64;
r2_68 <= r2_64;
r4_68 <= r4_64;
r5_68 <= r5_64;
r6_68 <= r6_64;
r7_68 <= r7_64;
r8_68 <= r8_64;
r9_68 <= r9_64;
r10_68 <= r10_64;
r11_68 <= r11_64;
r12_68 <= r12_64;
r13_68 <= r13_64;
r3_6c <= std_logic_vector( unsigned(r3_68) - unsigned(r1_68));
r0_6c <= r0_68;
r1_6c <= r1_68;
r2_6c <= r2_68;
r4_6c <= r4_68;
r5_6c <= r5_68;
r6_6c <= r6_68;
r7_6c <= r7_68;
r8_6c <= r8_68;
r9_6c <= r9_68;
r10_6c <= r10_68;
r11_6c <= r11_68;
r12_6c <= r12_68;
r13_6c <= r13_68;
r3_70 <= std_logic_vector(RESIZE(unsigned(r3_6c) * unsigned(r0_6c) + unsigned(r1_6c), 32));
r0_70 <= r0_6c;
r1_70 <= r1_6c;
r2_70 <= r2_6c;
r4_70 <= r4_6c;
r5_70 <= r5_6c;
r6_70 <= r6_6c;
r7_70 <= r7_6c;
r8_70 <= r8_6c;
r9_70 <= r9_6c;
r10_70 <= r10_6c;
r11_70 <= r11_6c;
r12_70 <= r12_6c;
r13_70 <= r13_6c;
t_70_s <= std_logic_vector(unsigned(r3_70) sll TO_INTEGER(unsigned(r0_70)));
r3_74 <= std_logic_vector( unsigned(r1_70) or unsigned(t_70_s));
r0_74 <= r0_70;
r1_74 <= r1_70;
r2_74 <= r2_70;
r4_74 <= r4_70;
r5_74 <= r5_70;
r6_74 <= r6_70;
r7_74 <= r7_70;
r8_74 <= r8_70;
r9_74 <= r9_70;
r10_74 <= r10_70;
r11_74 <= r11_70;
r12_74 <= r12_70;
r13_74 <= r13_70;
r3_78 <= std_logic_vector( unsigned(r3_74) xor unsigned(r0_74));
r0_78 <= r0_74;
r1_78 <= r1_74;
r2_78 <= r2_74;
r4_78 <= r4_74;
r5_78 <= r5_74;
r6_78 <= r6_74;
r7_78 <= r7_74;
r8_78 <= r8_74;
r9_78 <= r9_74;
r10_78 <= r10_74;
r11_78 <= r11_74;
r12_78 <= r12_74;
r13_78 <= r13_74;
r3_7c <= std_logic_vector( unsigned(r3_78) - unsigned(r1_78));
r0_7c <= r0_78;
r1_7c <= r1_78;
r2_7c <= r2_78;
r4_7c <= r4_78;
r5_7c <= r5_78;
r6_7c <= r6_78;
r7_7c <= r7_78;
r8_7c <= r8_78;
r9_7c <= r9_78;
r10_7c <= r10_78;
r11_7c <= r11_78;
r12_7c <= r12_78;
r13_7c <= r13_78;
r3_80 <= std_logic_vector(RESIZE(unsigned(r3_7c) * unsigned(r0_7c) + unsigned(r1_7c), 32));
r0_80 <= r0_7c;
r1_80 <= r1_7c;
r2_80 <= r2_7c;
r4_80 <= r4_7c;
r5_80 <= r5_7c;
r6_80 <= r6_7c;
r7_80 <= r7_7c;
r8_80 <= r8_7c;
r9_80 <= r9_7c;
r10_80 <= r10_7c;
r11_80 <= r11_7c;
r12_80 <= r12_7c;
r13_80 <= r13_7c;
t_80_s <= std_logic_vector(unsigned(r3_80) sll TO_INTEGER(unsigned(r0_80)));
r3_84 <= std_logic_vector( unsigned(r1_80) or unsigned(t_80_s));
r0_84 <= r0_80;
r1_84 <= r1_80;
r2_84 <= r2_80;
r4_84 <= r4_80;
r5_84 <= r5_80;
r6_84 <= r6_80;
r7_84 <= r7_80;
r8_84 <= r8_80;
r9_84 <= r9_80;
r10_84 <= r10_80;
r11_84 <= r11_80;
r12_84 <= r12_80;
r13_84 <= r13_80;
r3_88 <= std_logic_vector( unsigned(r3_84) xor unsigned(r0_84));
r0_88 <= r0_84;
r1_88 <= r1_84;
r2_88 <= r2_84;
r4_88 <= r4_84;
r5_88 <= r5_84;
r6_88 <= r6_84;
r7_88 <= r7_84;
r8_88 <= r8_84;
r9_88 <= r9_84;
r10_88 <= r10_84;
r11_88 <= r11_84;
r12_88 <= r12_84;
r13_88 <= r13_84;
r3_8c <= std_logic_vector( unsigned(r3_88) - unsigned(r1_88));
r0_8c <= r0_88;
r1_8c <= r1_88;
r2_8c <= r2_88;
r4_8c <= r4_88;
r5_8c <= r5_88;
r6_8c <= r6_88;
r7_8c <= r7_88;
r8_8c <= r8_88;
r9_8c <= r9_88;
r10_8c <= r10_88;
r11_8c <= r11_88;
r12_8c <= r12_88;
r13_8c <= r13_88;
r3_90 <= std_logic_vector(RESIZE(unsigned(r3_8c) * unsigned(r0_8c) + unsigned(r1_8c), 32));
r0_90 <= r0_8c;
r1_90 <= r1_8c;
r2_90 <= r2_8c;
r4_90 <= r4_8c;
r5_90 <= r5_8c;
r6_90 <= r6_8c;
r7_90 <= r7_8c;
r8_90 <= r8_8c;
r9_90 <= r9_8c;
r10_90 <= r10_8c;
r11_90 <= r11_8c;
r12_90 <= r12_8c;
r13_90 <= r13_8c;
t_90_s <= std_logic_vector(unsigned(r3_90) sll TO_INTEGER(unsigned(r0_90)));
r3_94 <= std_logic_vector( unsigned(r1_90) or unsigned(t_90_s));
r0_94 <= r0_90;
r1_94 <= r1_90;
r2_94 <= r2_90;
r4_94 <= r4_90;
r5_94 <= r5_90;
r6_94 <= r6_90;
r7_94 <= r7_90;
r8_94 <= r8_90;
r9_94 <= r9_90;
r10_94 <= r10_90;
r11_94 <= r11_90;
r12_94 <= r12_90;
r13_94 <= r13_90;
r3_98 <= std_logic_vector( unsigned(r3_94) xor unsigned(r0_94));
r0_98 <= r0_94;
r1_98 <= r1_94;
r2_98 <= r2_94;
r4_98 <= r4_94;
r5_98 <= r5_94;
r6_98 <= r6_94;
r7_98 <= r7_94;
r8_98 <= r8_94;
r9_98 <= r9_94;
r10_98 <= r10_94;
r11_98 <= r11_94;
r12_98 <= r12_94;
r13_98 <= r13_94;
r3_9c <= std_logic_vector( unsigned(r3_98) - unsigned(r1_98));
r0_9c <= r0_98;
r1_9c <= r1_98;
r2_9c <= r2_98;
r4_9c <= r4_98;
r5_9c <= r5_98;
r6_9c <= r6_98;
r7_9c <= r7_98;
r8_9c <= r8_98;
r9_9c <= r9_98;
r10_9c <= r10_98;
r11_9c <= r11_98;
r12_9c <= r12_98;
r13_9c <= r13_98;
r3_a0 <= std_logic_vector(RESIZE(unsigned(r3_9c) * unsigned(r0_9c) + unsigned(r1_9c), 32));
r0_a0 <= r0_9c;
r1_a0 <= r1_9c;
r2_a0 <= r2_9c;
r4_a0 <= r4_9c;
r5_a0 <= r5_9c;
r6_a0 <= r6_9c;
r7_a0 <= r7_9c;
r8_a0 <= r8_9c;
r9_a0 <= r9_9c;
r10_a0 <= r10_9c;
r11_a0 <= r11_9c;
r12_a0 <= r12_9c;
r13_a0 <= r13_9c;
t_a0_s <= std_logic_vector(unsigned(r3_a0) sll TO_INTEGER(unsigned(r0_a0)));
r3_a4 <= std_logic_vector( unsigned(r1_a0) or unsigned(t_a0_s));
r0_a4 <= r0_a0;
r1_a4 <= r1_a0;
r2_a4 <= r2_a0;
r4_a4 <= r4_a0;
r5_a4 <= r5_a0;
r6_a4 <= r6_a0;
r7_a4 <= r7_a0;
r8_a4 <= r8_a0;
r9_a4 <= r9_a0;
r10_a4 <= r10_a0;
r11_a4 <= r11_a0;
r12_a4 <= r12_a0;
r13_a4 <= r13_a0;
r3_a8 <= std_logic_vector( unsigned(r3_a4) xor unsigned(r0_a4));
r0_a8 <= r0_a4;
r1_a8 <= r1_a4;
r2_a8 <= r2_a4;
r4_a8 <= r4_a4;
r5_a8 <= r5_a4;
r6_a8 <= r6_a4;
r7_a8 <= r7_a4;
r8_a8 <= r8_a4;
r9_a8 <= r9_a4;
r10_a8 <= r10_a4;
r11_a8 <= r11_a4;
r12_a8 <= r12_a4;
r13_a8 <= r13_a4;
r3_ac <= std_logic_vector( unsigned(r3_a8) - unsigned(r1_a8));
r0_ac <= r0_a8;
r1_ac <= r1_a8;
r2_ac <= r2_a8;
r4_ac <= r4_a8;
r5_ac <= r5_a8;
r6_ac <= r6_a8;
r7_ac <= r7_a8;
r8_ac <= r8_a8;
r9_ac <= r9_a8;
r10_ac <= r10_a8;
r11_ac <= r11_a8;
r12_ac <= r12_a8;
r13_ac <= r13_a8;
r3_b0 <= std_logic_vector(RESIZE(unsigned(r3_ac) * unsigned(r0_ac) + unsigned(r1_ac), 32));
r0_b0 <= r0_ac;
r1_b0 <= r1_ac;
r2_b0 <= r2_ac;
r4_b0 <= r4_ac;
r5_b0 <= r5_ac;
r6_b0 <= r6_ac;
r7_b0 <= r7_ac;
r8_b0 <= r8_ac;
r9_b0 <= r9_ac;
r10_b0 <= r10_ac;
r11_b0 <= r11_ac;
r12_b0 <= r12_ac;
r13_b0 <= r13_ac;
t_b0_s <= std_logic_vector(unsigned(r3_b0) sll TO_INTEGER(unsigned(r0_b0)));
r3_b4 <= std_logic_vector( unsigned(r1_b0) or unsigned(t_b0_s));
r0_b4 <= r0_b0;
r1_b4 <= r1_b0;
r2_b4 <= r2_b0;
r4_b4 <= r4_b0;
r5_b4 <= r5_b0;
r6_b4 <= r6_b0;
r7_b4 <= r7_b0;
r8_b4 <= r8_b0;
r9_b4 <= r9_b0;
r10_b4 <= r10_b0;
r11_b4 <= r11_b0;
r12_b4 <= r12_b0;
r13_b4 <= r13_b0;
r3_b8 <= std_logic_vector( unsigned(r3_b4) xor unsigned(r0_b4));
r0_b8 <= r0_b4;
r1_b8 <= r1_b4;
r2_b8 <= r2_b4;
r4_b8 <= r4_b4;
r5_b8 <= r5_b4;
r6_b8 <= r6_b4;
r7_b8 <= r7_b4;
r8_b8 <= r8_b4;
r9_b8 <= r9_b4;
r10_b8 <= r10_b4;
r11_b8 <= r11_b4;
r12_b8 <= r12_b4;
r13_b8 <= r13_b4;
r3_bc <= std_logic_vector( unsigned(r3_b8) - unsigned(r1_b8));
r0_bc <= r0_b8;
r1_bc <= r1_b8;
r2_bc <= r2_b8;
r4_bc <= r4_b8;
r5_bc <= r5_b8;
r6_bc <= r6_b8;
r7_bc <= r7_b8;
r8_bc <= r8_b8;
r9_bc <= r9_b8;
r10_bc <= r10_b8;
r11_bc <= r11_b8;
r12_bc <= r12_b8;
r13_bc <= r13_b8;
r3_c0 <= std_logic_vector(RESIZE(unsigned(r3_bc) * unsigned(r0_bc) + unsigned(r1_bc), 32));
r0_c0 <= r0_bc;
r1_c0 <= r1_bc;
r2_c0 <= r2_bc;
r4_c0 <= r4_bc;
r5_c0 <= r5_bc;
r6_c0 <= r6_bc;
r7_c0 <= r7_bc;
r8_c0 <= r8_bc;
r9_c0 <= r9_bc;
r10_c0 <= r10_bc;
r11_c0 <= r11_bc;
r12_c0 <= r12_bc;
r13_c0 <= r13_bc;
t_c0_s <= std_logic_vector(unsigned(r3_c0) sll TO_INTEGER(unsigned(r0_c0)));
r3_c4 <= std_logic_vector( unsigned(r1_c0) or unsigned(t_c0_s));
r0_c4 <= r0_c0;
r1_c4 <= r1_c0;
r2_c4 <= r2_c0;
r4_c4 <= r4_c0;
r5_c4 <= r5_c0;
r6_c4 <= r6_c0;
r7_c4 <= r7_c0;
r8_c4 <= r8_c0;
r9_c4 <= r9_c0;
r10_c4 <= r10_c0;
r11_c4 <= r11_c0;
r12_c4 <= r12_c0;
r13_c4 <= r13_c0;
r3_c8 <= std_logic_vector( unsigned(r3_c4) xor unsigned(r0_c4));
r0_c8 <= r0_c4;
r1_c8 <= r1_c4;
r2_c8 <= r2_c4;
r4_c8 <= r4_c4;
r5_c8 <= r5_c4;
r6_c8 <= r6_c4;
r7_c8 <= r7_c4;
r8_c8 <= r8_c4;
r9_c8 <= r9_c4;
r10_c8 <= r10_c4;
r11_c8 <= r11_c4;
r12_c8 <= r12_c4;
r13_c8 <= r13_c4;
r3_cc <= std_logic_vector( unsigned(r3_c8) - unsigned(r1_c8));
r0_cc <= r0_c8;
r1_cc <= r1_c8;
r2_cc <= r2_c8;
r4_cc <= r4_c8;
r5_cc <= r5_c8;
r6_cc <= r6_c8;
r7_cc <= r7_c8;
r8_cc <= r8_c8;
r9_cc <= r9_c8;
r10_cc <= r10_c8;
r11_cc <= r11_c8;
r12_cc <= r12_c8;
r13_cc <= r13_c8;
r3_d0 <= std_logic_vector(RESIZE(unsigned(r3_cc) * unsigned(r0_cc) + unsigned(r1_cc), 32));
r0_d0 <= r0_cc;
r1_d0 <= r1_cc;
r2_d0 <= r2_cc;
r4_d0 <= r4_cc;
r5_d0 <= r5_cc;
r6_d0 <= r6_cc;
r7_d0 <= r7_cc;
r8_d0 <= r8_cc;
r9_d0 <= r9_cc;
r10_d0 <= r10_cc;
r11_d0 <= r11_cc;
r12_d0 <= r12_cc;
r13_d0 <= r13_cc;
t_d0_s <= std_logic_vector(unsigned(r3_d0) sll TO_INTEGER(unsigned(r0_d0)));
r3_d4 <= std_logic_vector( unsigned(r1_d0) or unsigned(t_d0_s));
r0_d4 <= r0_d0;
r1_d4 <= r1_d0;
r2_d4 <= r2_d0;
r4_d4 <= r4_d0;
r5_d4 <= r5_d0;
r6_d4 <= r6_d0;
r7_d4 <= r7_d0;
r8_d4 <= r8_d0;
r9_d4 <= r9_d0;
r10_d4 <= r10_d0;
r11_d4 <= r11_d0;
r12_d4 <= r12_d0;
r13_d4 <= r13_d0;
r0_d8 <= std_logic_vector( unsigned(r0_d4) xor unsigned(r3_d4));
r1_d8 <= r1_d4;
r2_d8 <= r2_d4;
r3_d8 <= r3_d4;
r4_d8 <= r4_d4;
r5_d8 <= r5_d4;
r6_d8 <= r6_d4;
r7_d8 <= r7_d4;
r8_d8 <= r8_d4;
r9_d8 <= r9_d4;
r10_d8 <= r10_d4;
r11_d8 <= r11_d4;
r12_d8 <= r12_d4;
r13_d8 <= r13_d4;
r0_dc <= std_logic_vector( unsigned(r0_d8) - unsigned(r1_d8));
regs_out(0) <= r0_d8;
regs_out(1) <= r1_d8;
regs_out(2) <= r2_d8;
regs_out(3) <= r3_d8;
regs_out(4) <= r4_d8;
regs_out(5) <= r5_d8;
regs_out(6) <= r6_d8;
regs_out(7) <= r7_d8;
regs_out(8) <= r8_d8;
regs_out(9) <= r9_d8;
regs_out(10) <= r10_d8;
regs_out(11) <= r11_d8;
regs_out(12) <= r12_d8;
regs_out(13) <= r13_d8;

--->>> END LOGIC

end architecture offload_top_1;

